��  CCircuit��  CSerializeHack           ��  CPart    �   �     ���  CNAND�� 	 CTerminal  ����              @          
�  ��	              @          
�   !               �            ��           ��    �� 	 CLogicOut
�  �0�1               �            �(�8           ��    ��  CLogicIn�� 	 CLatchKey  xi�w         
�  �p�q                            �l�t         ����     ��  x!�/        
�  �(�)              @            �$�,        ����     ��  x���        
�  ����              @            ����        ����     ��  COR
�  h(})               �          
�  h8}9                          
�  �0�1               �            |$�<           ��        �   �     ���  CWire  �0�1      "�  h i)       "�    i      "�  h8iq       "�  �piq      "�  ��)       "�  �(�)      "�  ����          �   �     �    �   �         �   �      *   (    %  #    '   )   *  $   &      #    %   $  '  &  )  (               �$s�        @     +        @            @    "V  (      �                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 