��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CLogicOut�� 	 CTerminal  `XuY      	       @            tP�`          ��    ��  CLogicIn�� 	 CLatchKey  py��         
�  ����                            �|��         ����     ��  pa�o         
�  �h�i                            �d�l         ����     ��  pA�O         
�  �H�I                            �D�L         ����     ��  COR
�   P5Q      	       @          
�   `5a                          
�  LXaY              @            4LLd           ��    �� 	 CInverter
�  �H�I      	                   
�  �H�I              @            �<�T           ��    ��  CNAND
�  �H�I      	       @          
�  �X�Y                          
�  P!Q              @            �D\     "      ��                  ���  CWire   `!�       &�  ��!�      &�  �X�i       &�  �h�i                    �                                 (   *     $   '          " "  " # ) # $ $   (  ' # *  )             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 