��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CLogicOut�� 	 CTerminal  0$19              @            (8$         ��    ��  CLogicIn�� 	 CLatchKey  HQX_        
�  dXyY              @            \Td\        ����     ��  H�X�        
�  d�y�              @            \�d�        ����     ��  H	X        
�  dy              @            \d        ����     ��  CAND
�  @HUI              @          
�  @XUY               �          
�  lP�Q               �            TDl\           ��    ��  COR
�  ��              @          
�  � �!              @          
�                @            �$           ��    ��  CNAND
�  ����              @          
�  ����              @          
�  ��               �            ���     #      ��    �� 	 CInverter
�  �P�Q               �          
�  �PQ              @            �D�\     (      ��                  ���  CWire  081Q       +�   P1Q      +�  �P�Q      +�  XAY      +�  X�       +�  HAI      +�  I       +�  xX�Y      +�  � �Y       +�  ����       +�  x���      +�  �X��       +�  x�                    �                              ,   3   6   8  1   /    .  8   4      2 # 7 # $ 5 $ % % 0 ( . ( ) ) -  - ) ,  ( 0  / % 2    1  7  3 $ 6  5 4 #               �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 