��  CCircuit��  CSerializeHack           ��  CPart              ���  CAND�� 	 CTerminal   �5�              @          
�   �5�              @          
�  L�a�              @            4�L�           ��    �� 	 CLogicOut
�   PQ              @            H$X          ��    ��  CLogicIn�� 	 CLatchKey  `�p�        
�  |���              @            t�|�        ����     ��  `apo         
�  |h�i                            td|l         ����     �
�  �H�I              @          
�  �X�Y              @          
�  �P�Q              @            �D�\           ��    ��  `!p/         
�  |(�)                            t$|,         ����     ��  CNAND
�  �01                          
�  �@A                          
�  819              @            ,D     "      ��                  ���  CWire  �PQ      &�  `X�Y      &�  `Xa�       &�  0H�I      &�  081I       &�  ��!�      &�  ����      &�  ����       &�  ��!�      &�   �!�       &�  �@�i       &�  �h�i      &�  �(�1       &�  �(�)                    �                             0   /    )  '    -   2  *   (    '   4 " 3 " # 1 # $ $ +   )  (  +  $ * - 0  . , / .   , # 2  1 4 "  3             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 